`timescale 1 ns / 1 ps

module AESL_deadlock_detector (
    input reset,
    input clock);

    wire [0:0] proc_dep_vld_vec_0;
    reg [0:0] proc_dep_vld_vec_0_reg;
    wire [0:0] in_chan_dep_vld_vec_0;
    wire [1:0] in_chan_dep_data_vec_0;
    wire [0:0] token_in_vec_0;
    wire [0:0] out_chan_dep_vld_vec_0;
    wire [1:0] out_chan_dep_data_0;
    wire [0:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [1:0] dep_chan_data_1_0;
    wire token_1_0;
    wire [0:0] proc_dep_vld_vec_1;
    reg [0:0] proc_dep_vld_vec_1_reg;
    wire [0:0] in_chan_dep_vld_vec_1;
    wire [1:0] in_chan_dep_data_vec_1;
    wire [0:0] token_in_vec_1;
    wire [0:0] out_chan_dep_vld_vec_1;
    wire [1:0] out_chan_dep_data_1;
    wire [0:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [1:0] dep_chan_data_0_1;
    wire token_0_1;
    wire [1:0] dl_in_vec;
    wire dl_detect_out;
    wire [1:0] origin;
    wire token_clear;

    reg ap_done_reg_0;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_0 <= 'b0;
        end
        else begin
            ap_done_reg_0 <= AESL_inst_myFuncAccel.Block_codeRepl93_pro_U0.ap_done;
        end
    end

    reg ap_done_reg_1;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_1 <= 'b0;
        end
        else begin
            ap_done_reg_1 <= AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_done;
        end
    end

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myFuncAccel$Block_codeRepl93_pro_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myFuncAccel$Block_codeRepl93_pro_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myFuncAccel$Block_codeRepl93_pro_U0$ap_idle <= AESL_inst_myFuncAccel.Block_codeRepl93_pro_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myFuncAccel.Block_codeRepl93_pro_U0
    AESL_deadlock_detect_unit #(2, 0, 1, 1) AESL_deadlock_detect_unit_0 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (~AESL_inst_myFuncAccel.empty_U.i_full_n & AESL_inst_myFuncAccel.Block_codeRepl93_pro_U0.ap_done & deadlock_detector.ap_done_reg_0 & ~AESL_inst_myFuncAccel.empty_U.t_read | ((AESL_inst_myFuncAccel.Block_codeRepl93_pro_U0_ap_ready_count[0]) & AESL_inst_myFuncAccel.Block_codeRepl93_pro_U0.ap_idle & ~(AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0_ap_ready_count[0])));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[1 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[0];

    // delay ap_idle for one cycle
    reg [0:0] AESL_inst_myFuncAccel$Loop_sizeLoop_proc_U0$ap_idle;
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            AESL_inst_myFuncAccel$Loop_sizeLoop_proc_U0$ap_idle <= 'b0;
        end
        else begin
            AESL_inst_myFuncAccel$Loop_sizeLoop_proc_U0$ap_idle <= AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle;
        end
    end
    // Process: AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0
    AESL_deadlock_detect_unit #(2, 1, 1, 1) AESL_deadlock_detect_unit_1 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (~AESL_inst_myFuncAccel.empty_U.t_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.empty_U.i_write | ~AESL_inst_myFuncAccel.data0_load_6_loc_cha_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_6_loc_cha_U.if_write | ~AESL_inst_myFuncAccel.data0_load_7_loc_cha_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_7_loc_cha_U.if_write | ~AESL_inst_myFuncAccel.data0_load_8_loc_cha_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_8_loc_cha_U.if_write | ~AESL_inst_myFuncAccel.data0_load_9_loc_cha_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_9_loc_cha_U.if_write | ~AESL_inst_myFuncAccel.data0_load_10_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_10_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_11_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_11_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_12_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_12_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_13_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_13_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_14_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_14_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_15_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_15_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_16_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_16_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_17_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_17_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_18_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_18_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_19_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_19_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_20_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_20_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_21_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_21_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_22_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_22_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_23_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_23_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_24_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_24_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_25_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_25_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_26_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_26_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_27_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_27_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_28_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_28_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_29_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_29_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_30_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_30_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_31_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_31_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_32_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_32_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_33_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_33_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_34_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_34_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_35_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_35_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_36_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_36_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_37_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_37_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_38_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_38_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_39_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_39_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_40_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_40_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_41_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_41_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_42_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_42_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_43_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_43_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_44_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_44_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_45_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_45_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_46_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_46_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_47_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_47_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_48_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_48_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_49_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_49_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_50_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_50_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_51_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_51_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_52_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_52_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_53_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_53_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_54_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_54_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_55_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_55_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_56_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_56_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_57_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_57_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_58_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_58_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_59_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_59_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_60_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_60_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_61_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_61_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_62_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_62_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_63_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_63_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_64_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_64_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_65_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_65_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_66_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_66_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_67_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_67_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_68_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_68_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_69_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_69_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_70_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_70_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_71_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_71_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_72_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_72_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_73_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_73_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_74_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_74_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_75_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_75_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_76_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_76_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_77_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_77_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_78_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_78_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_79_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_79_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_80_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_80_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_81_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_81_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_82_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_82_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_83_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_83_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_84_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_84_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_85_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_85_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_86_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_86_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_87_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_87_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_88_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_88_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_89_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_89_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_90_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_90_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_91_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_91_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_92_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_92_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_93_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_93_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_94_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_94_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_95_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_95_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_96_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_96_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_97_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_97_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_98_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_98_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_99_loc_ch_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_99_loc_ch_U.if_write | ~AESL_inst_myFuncAccel.data0_load_100_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_100_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_101_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_101_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_102_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_102_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_103_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_103_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_104_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_104_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_105_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_105_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_106_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_106_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_107_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_107_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_108_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_108_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_109_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_109_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_110_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_110_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_111_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_111_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_112_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_112_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_113_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_113_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_114_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_114_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_115_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_115_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_116_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_116_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_117_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_117_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_118_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_118_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_119_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_119_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_120_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_120_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_121_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_121_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_122_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_122_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_123_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_123_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_124_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_124_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_125_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_125_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_126_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_126_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_127_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_127_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_128_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_128_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_129_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_129_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_130_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_130_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_131_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_131_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_132_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_132_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_133_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_133_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_134_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_134_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_135_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_135_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_136_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_136_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_137_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_137_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_138_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_138_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_139_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_139_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_140_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_140_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_141_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_141_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_142_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_142_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_143_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_143_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_144_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_144_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_145_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_145_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_146_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_146_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_147_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_147_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_148_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_148_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_149_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_149_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_150_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_150_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_151_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_151_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_152_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_152_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_153_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_153_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_154_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_154_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_155_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_155_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_156_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_156_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_157_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_157_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_158_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_158_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_159_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_159_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_160_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_160_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_161_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_161_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_162_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_162_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_163_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_163_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_164_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_164_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_165_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_165_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_166_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_166_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_167_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_167_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_168_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_168_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_169_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_169_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_170_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_170_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_171_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_171_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_172_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_172_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_173_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_173_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_174_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_174_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_175_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_175_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_176_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_176_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_177_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_177_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_178_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_178_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_179_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_179_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_180_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_180_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_181_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_181_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_182_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_182_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_183_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_183_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_184_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_184_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_185_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_185_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_186_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_186_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_187_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_187_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_188_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_188_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_189_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_189_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_190_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_190_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_191_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_191_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_192_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_192_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_193_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_193_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_194_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_194_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_195_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_195_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_196_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_196_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_197_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_197_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_198_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_198_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_199_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_199_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_200_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_200_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_201_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_201_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_202_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_202_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_203_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_203_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_204_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_204_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_205_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_205_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_206_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_206_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_207_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_207_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_208_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_208_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_209_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_209_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_210_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_210_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_211_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_211_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_212_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_212_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_213_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_213_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_214_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_214_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_215_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_215_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_216_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_216_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_217_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_217_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_218_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_218_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_219_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_219_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_220_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_220_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_221_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_221_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_222_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_222_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_223_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_223_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_224_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_224_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_225_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_225_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_226_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_226_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_227_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_227_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_228_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_228_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_229_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_229_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_230_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_230_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_231_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_231_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_232_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_232_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_233_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_233_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_234_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_234_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_235_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_235_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_236_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_236_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_237_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_237_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_238_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_238_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_239_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_239_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_240_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_240_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_241_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_241_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_242_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_242_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_243_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_243_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_244_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_244_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_245_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_245_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_246_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_246_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_247_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_247_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_248_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_248_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_249_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_249_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_250_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_250_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_251_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_251_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_252_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_252_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_253_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_253_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_254_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_254_loc_c_U.if_write | ~AESL_inst_myFuncAccel.data0_load_255_loc_c_U.if_empty_n & (AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_ready | AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle) & ~AESL_inst_myFuncAccel.data0_load_255_loc_c_U.if_write | ((AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0_ap_ready_count[0]) & AESL_inst_myFuncAccel.Loop_sizeLoop_proc_U0.ap_idle & ~(AESL_inst_myFuncAccel.Block_codeRepl93_pro_U0_ap_ready_count[0])));
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[1 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[0];


    AESL_deadlock_report_unit #(2) AESL_deadlock_report_unit_inst (
        .reset(reset),
        .clock(clock),
        .dl_in_vec(dl_in_vec),
        .dl_detect_out(dl_detect_out),
        .origin(origin),
        .token_clear(token_clear));

endmodule
